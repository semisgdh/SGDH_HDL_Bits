module top_module (
    output zero  // 출력 신호 선언
);
    assign zero = 1'b0;  // 항상 0을 출력
endmodule